* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Inductors
L1 1 2 
L2 2 4 2.1529p
L3 4 6 1.9729p
L4 6 8 2.3966p
L5 8 10 1.6354p
L6 13 14 2.2793p
L7 15 16
L8 16 18 2.1529p
L9 18 20 1.9729p
L10 20 22 2.3966p
L11 22 24 1.6354p
L12 27 14 2.2793p
L13 31 32
L14 32 34 2.2381p
L15 34 36 2.0205p
L16 36 38 2.0178p
L17 38 40 1.8033p
L18 43 30 2.2246p
L19 14 29 1.7515p
L20 30 45 3.8658p
L21 45 48 
LP1 3 0
LP2 7 0
LP3 9 0
LP4 11 0
LP6 17 0
LP7 21 0
LP8 23 0
LP9 25 0
LP11 33 0
LP12 37 0
LP13 39 0
LP14 41 0
LP17 44 0
LP18 46 0
LB1 4 5
LB2 10 12
LB3 18 19
LB4 24 26
LB5 34 35
LB6 40 42
LB7 14 28
LB8 45 47
* Ports
P1 1 0
P2 15 0
P3 31 0
P4 48 0
PB1 5 0
PB2 12 0
PB3 19 0
PB4 26 0
PB5 35 0
PB6 42 0
PB7 28 0
PB8 47 0
J1 2 3 121u
J2 6 7 116u
J3 8 9 90u
J4 10 11 280u
J5 10 13 192u
J6 16 17 121u
J7 20 21 116u
J8 22 23 90u
J9 24 25 280u
J10 24 27 192u
J11 32 33 72u
J12 36 37 77u
J13 38 39 83u
J14 40 41 169u
J15 40 43 129u
J16 29 30 149u
J17 30 44 93u
J18 45 46 137u
.end