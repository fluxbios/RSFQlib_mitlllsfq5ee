* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Inductors
L1 1 2
L2 2 4 4.0481p
L3 4 6 3.6036p
L4 6 8 7.2183p
L5 8 11 3.0677p
L7 12 29 2.5596p
L8 16 17 
L9 17 19 4.0481p
L10 19 21 3.6036p
L11 21 23 4.3879p
L12 23 26 3.217p
L13 27 29 3.2439p
L14 33 34 
L15 34 36 4.3135p
L16 36 38 3.926p
L17 38 40 7.5833p
L18 40 42 1.2875p
L19 42 44 1.0678p
L21 30 31 0.37382p
L22 31 46 0.52995p
L23 46 47 0.95137p
L24 47 49 2.5089p
L25 49 51 1.2791p
L26 51 53 3.5427p
L27 53 56 
LP1 3 0
LP2 7 0
LP3 9 0
LP5 13 0
LP6 18 0
LP7 22 0
LP8 24 0
LP10 28 0
LP12 35 0
LP13 39 0
LP14 41 0
LP16 48 0
LP17 52 0
LP18 54 0
LB1 4 5
LB2 8 10
LB3 12 15
LB4 19 20
LB5 23 25
LB6 36 37
LB7 42 43
LB8 31 32
LB9 49 50
LB10 53 55

* Ports
P1 1 0
P2 16 0
P3 33 0
P4 56 0
PB1 5 0
PB2 10 0
PB3 15 0
PB4 20 0
PB5 25 0
PB6 37 0
PB7 43 0
PB8 32 0
PB9 50 0
PB10 55 0
J1 2 3 86u
J2 6 7 100u
J3 8 9 191u
J4 11 12 178u
J5 12 13 116u
J6 17 18 86u
J7 21 22 100u
J8 23 24 235u
J9 26 27 196u
J10 27 28 284u
J11 29 30 78u
J12 34 35 99u
J13 38 39 94u
J14 40 41 218u
J15 44 46 165u
J16 47 48 163u
J17 51 52 151u
J18 53 54 236u
.end