* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Inductors
L1 1 2 
L2 2 6 5.2p
L3 6 9 2.07p 
L4 9 11 2.07p
L5 11 14
LB1 2 5 
LB2 9 10 
LP1 3 0 
LP2 7 0 
LP3 12 0 
* Ports
P1 1 0
P2 14 0
PB1 5 0
PB2 10 0
J1 2 3 200u
J2 6 7 250u
J3 11 12 250u
.end