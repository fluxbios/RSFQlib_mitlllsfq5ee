* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Inductors
L1 1 2 2p
L2 2 4 2p	
L3 4 6 1p	
L4 6 7 2.3p
L5 7 9 2p	
L6 6 10 2.3p
L7 10 12 2p	
LP1 3 0
LP2 8 0
LP3 11 0
LB1 4 5
* Ports
P1 1 0
P2 9 0
P3 12 0
PB1 5 0
J1 2 3 325u
J2 7 8 150u
J3 10 11 150u
.end