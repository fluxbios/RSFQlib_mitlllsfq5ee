* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Inductors
L1 1 2 2.5p
L2 2 5 3.3p
L3 5 8 
LP1 3 0
LP2 6 0
LB1 2 4
LB2 5 7
* Ports
P1 1 0
P2 4 0
P3 7 0
P4 8 0
J1 2 3	200u
J2 5 6	162u
.end