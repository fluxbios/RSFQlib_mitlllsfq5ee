* Circuit for InductEx extraction (excluding resistors)
* Author: L. Schindler
* Version: 1.5.1
* Last modification date: 18 June 2020
* Last modification by: L. Schindler

* Inductors
L1 1 2				
L2 2 4 2.0822p		
L3 4 6 2.6809p		
L4 8 9 1.3486p		
L5 10 11			
L6 11 13 2.0822p	
L7 13 15 2.6809p	
L8 43 9 1.3486p		
L10 9 19 1.8890p	
L12 22 24 5.4916p	
L13 25 26		
L14 26 28 3.3652p
L15 28 30 4.0267p	
L16 30 32			
L17 24 33 1.5727p	
L18 33 35 2.0776p	
L19 35 37 0.885p	
L20 37 39 4.2904p
L21 39 42			
LB1 4 5			
LB2 13 14		
LB3 9 18			
LB4 22 23			
LB5 28 29			
LB6 35 36			
LB7 39 40			
LP1 3 0			
LP2 7 0				
LP4 12 0			
LP5 16 0			
LP8 21 0		
LP9 27 0		
LP10 31 0			
LP12 34 0			
LP13 38 0			
LP14 41 0			
* Ports
P1 1 0
P2 10 0
P3 25 0
P4 42 0
PB1 5 0
PB2 14 0
PB3 18 0
PB4 23 0
PB5 29 0
PB6 36 0
PB7 40 0
J1 2 3  	117u
J2 6 7  	195u
J3 6 8		131u
J4 11 12	117u
J5 15 16	195u
J6 15 43	131u
J7 19 22	220u
J8 22 21	172u
J9 26 27	081u
J10 30 31	075u
J11 32 24	063u
J12 33 34	140u
J13 37 38	162u
J14 39 41	190u
.end